module pfd (input ref_clk, input gated_dco_clk, input sample, output early,output early_edge, output late_edge);
endmodule // pfd
